module model_config_mem
(
    input clk_i,
    input rst_ni,


);

endmodule